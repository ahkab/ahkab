TEST
vs 1 0 type=sin 0 15 60 0 0 
rload 1 0 10k
.tran tstep=1m tstop=30m 
*.plot tran v(1) 
.fft I(VS) np=512
.end
