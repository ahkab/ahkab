* Cockcroft-Walton x8 multiplier
D1 7 8 d
C1 8 6 1000p
D2 6 7 d
C2 5 7 1000p
D3 5 6 d
C3 4 6 1000p
D4 4 5 d
C4 3 5 1000p
D5 3 4 d
C5 2 4 1000p
D6 2 3 d
D7 1 2 d
C6 1 3 1000p
C7 2 0 1000p
C8 99 1 1000p
D8 0 1 d
V1 99 0 type=vdc vdc=0 type=SIN vo=0 va=5 freq=1k
.model diode d
.op
.tran 0.01m 50m
.plot tran v(8) v(6) v(4) v(2)
.end
