Untitled
R0 n2 0 820000
C1 n3 0 3.9e-11
R1 n3 n1 51000000
R2 n1 n4 220000
R3 0 n4 6200000
R4 n4 n3 13000
L1 n6 0 1.3e-08
C2 n3 n4 3.9e-07
V1 n1 0 type=vdc vdc=5 vac=1 type=pulse v1=0 v2=1 td=5e-07 per=2 tr=1e-12 tf=1e-12 pw=1

.op
.ac start=1e3 stop=1e5 nsteps=10