Untitled
L0 0 n4 4e-09
L1 0 n3 3.6e-08
R0 0 n1 10
C0 n4 n1 1.5e-10
L2 n1 n3 1.5e-08
R1 n2 0 390
L3 0 0 7e-09
V1 n1 0 type=vdc vdc=5 vac=1 type=pulse v1=0 v2=1 td=5e-07 per=2 tr=1e-12 tf=1e-12 pw=1

.op
.ac start=1e3 stop=1e5 nsteps=10