** PZ TEST
IN   0  1  type=idc idc=1.00  iac=1
R1   1  0  1.0
C3   1  0  1.52
C4   2  0  1.50
C5   3  0  0.83
C1   1  2  0.93
L1   1  2  0.65
C2   2  3  3.80
L2   2  3  1.00
R2   3  4  1.00
VT   4  0  type=vdc vdc=0
.PZ  V(4,0) IN
*.AC  DEC  100  .001HZ  10HZ
*.PLOT AC  IDB(R2)  IP(R2)
.END
 
