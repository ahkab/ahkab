MOS COLPITTS OSCILLATOR

vdd dd 0 type=vdc vdc=2.5

* Ql = 33 at 3GHz
L1 dd nd 5n ic=-1n
R0 nd dd 3.5k 

* n = 0.5, f0 = 3GHz
C1 nd ns 1.12p ic=2.5
C2 ns 0  1.12p *ic=.01

m1 nd1 bias ns ns nmos w=200u l=1u
vtest nd nd1 type=vdc vdc=0 *read current

* Bias
vbias bias 0 type=vdc vdc=2
ib ns 0 type=idc idc=1.3m

.model ekv nmos TYPE=n VTO=.4 KP=10e-6

.op
.tran tstop=250n tstep=.1n method=trap uic=2
*.plot tran v(nd)
