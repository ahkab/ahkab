RC time delay circuit
v1 1 0 type=vdc vdc=0 type=pulse v1=0 v2=10 td=0 tr=10n tf=1p pw=100 per=1000
c1 2 0 55p ic=0
*c2 1 2 22u ic=0
r1 2 1 33k
.op
.tran tstep=100n tstop=10u uic=2
.plot tran v(2) v(1,2)
*.print tran v(1,2)
.end 

