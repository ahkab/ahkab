** PZ TEST
IN   0  1  type=idc idc=1.00  iac=1
R1   1  0  1.0
C3   1  0  1.52
C4   2  0  1.50
C5   3  0  0.83
C1   1  2  0.93
L1   1  2  0.65
C2   2  3  3.80
L2   2  3  1.00
R2   3  0  1.00
.PZ  V(3,0) IN
.AC nsteps=100 start=.1 stop=10
.plot ac |v(3)|
.END
 
