FILE: FLP9TH.SP
******

VIN  IN  0  AC 1
.PZ  V(OUT) VIN
.AC  DEC  50  .1K  100K
.OPTIONS  POST  DCSTEP=1E3  X0R=-1.23456E+3  X1R=-1.23456E+2
+ X2R=1.23456E+3  FSCAL=1E-6  GSCAL=1E3  CSCAL=1E9  LSCAL=1E3
.PLOT  AC  VDB(OUT)

.SUBCKT OPAMP IN+ IN- OUT GM1=2 RI=1K CI=26.6U GM2=1.33333 RL=75
RII IN+ IN- 2MEG
RI1 IN+ 0 500MEG
RI2 IN- 0 500MEG
G1  1  0  IN+  IN-  GM1
C1  1  0  CI
R1  1  0  RI
G2   OUT  0  1  0  GM2
RLD  OUT  0  RL
.ENDS

.SUBCKT FDNR 1 R1=2K C1=12N R4=4.5K 
RLX=75
R1  1  2  R1
C1  2  3  C1
R2  3  4  3.3K
R3  4  5  3.3K
R4  5  6  R4
C2  6  0  10N
XOP1  2  4  5  OPAMP
XOP2  6  4  3  OPAMP
.ENDS

*

RS IN 1 5.4779K
R12 1 2 4.44K
R23 2 3 3.2201K
R34 3 4 3.63678K
R45 4 OUT 1.2201K
C5 OUT 0 10N

X1 1 FDNR R1=2.0076K  C1=12N    R4=4.5898K
X2 2 FDNR R1=5.9999K  C1=6.8N   R4=4.25725K
X3 3 FDNR R1=5.88327K C1=4.7N   R4=5.62599K
X4 4 FDNR R1=1.0301K  C1=6.8N   R4=5.808498K

.END


