* Shooting solution

.include diffamp.spc

.op
