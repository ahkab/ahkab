KERWIN'S CIRCUIT HAVING JW-AXIS TRANSMISSION ZEROS.

**
* T = V(5) / VIN
*   = 1.2146 (S**2 + 2) / (S**2 + 0.1*S + 1)
* POLES = (-0.05004, +0.9987), (-0.05004, -0.9987)
* ZEROS = (0.0, +1.4142), (0.0, -1.4142)
*****

VIN  1  0  type=vdc vdc=1
C1   1  2  0.7071
C2   2  4  0.7071
C3   3  0  1.4142 
C4   4  0  0.3536
R1   1  3  1.0
R2   3  4  1.0
R3   2  5  0.5
E1   5  0  4  0  2.4293
.OP
.PZ  V(5,0)  VIN
.END
