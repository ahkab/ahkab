5TH-ORDER LOW_PASS FILTER
****
* T = I(R2) / IIN
*   = 0.113*(S**2 + 1.6543)*(S**2 + 0.2632) /
*     (S**5 + 0.9206*S**4 + 1.26123*S**3 +
*      0.74556*S**2 + 0.2705*S  + 0.09836)
*****
IN   0  1  type=idc idc=1.00
R1   1  0  1.0
C3   1  0  1.52
C4   2  0  1.50
C5   3  0  0.83
C1   1  2  0.93
L1   1  2  0.65
C2   2  3  3.80
L2   2  3  1.00
R2   3  0  1.00
.OP
.PZ  V(3,0) IN
.END
