*FILE: FHP4TH.SP
*****
* T = V(10) / VIN
*  = (S**4) / ((S**2 + 0.7653*S + 1) * (S**2 + 1.8477*S + 1))
*
* POLES, (-0.38265, +0.923895), (-0.38265, -0.923895)
*          (-0.9239, +0.3827),   (-0.9239, -0.3827)
* ZEROS, FOUR ZEROS AT (0.0, 0.0)
*****

VIN  1  0  type=vdc vdc=1
C1   1  2  1
C2   2  3  1
R1   3  0  2.613
R2   2  4  0.3826
E1   4  0  3  0  1
C3   4  5  1
C4   5  6  1
R3   6  0  1.0825
R4   5  10 0.9238
E2   10 0  6  0  1
RL   10 0  1E20

.PZ   V(10,0)   VIN 
.END
